`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:04:26 09/23/2013 
// Design Name: 
// Module Name:    top_level 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top_level(
    input clk,
    input rst,
	 input  [7:0] p0,p1,p2,p3,p5,p6,p7,p8,
	 output [7:0] out_data

);

wire signed [10:0] gx, gy;    // 11 bit: gx es gy max ertekei: 255*4 + elojel
wire signed [10:0] abs_gx, abs_gy;	// absz.ertek
wire [10:0] sum;				  // kimenet: max 255*8 bit lehet

assign gx =((p2-p0) + ((p5-p3)<<1) + (p8-p6));		// sobel mask for gradient in horiz. direction
assign gy =((p0-p6) + ((p1-p7)<<1) + (p2-p8));		// sobel mask for gradient in vertical direction

assign abs_gx = (gx[10] ? ~gx+1 : gx);					// ha negativ: absz erteket veszem
assign abs_gy = (gy[10] ? ~gy+1 : gy);	

assign sum = abs_gx + abs_gy;							// x es y irany osszeadasa

assign out_data = (|sum[10:8]) ? 8'hff : sum[7:0];	// 255 lehet a max ertek

endmodule



/*reg [7:0] first_row [255:0];
reg [7:0] cntr;
always @ (posedge clk)
begin
	if(rst | cntr == 255)
		cntr <= 0;
	else 
		cntr <= cntr + 1;
end

reg [7:0] konv_input [2:0][2:0];

always @ (posedge clk)
begin
	
		first_row[cntr] <= data_in;
end*/

